r1 out 0 1
v1 in 0 100
n1 in 0 out 0 10

