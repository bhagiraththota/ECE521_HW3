vdd 1 0 5
r1 1 2 1000
d1 2 3 dmod 1
va 3 0 5
d2 2 0 dmod 1
d3 2 4 dmod 1
r2 4 0 1000
