vdd 1 0 5
mp1 2 3 1 1 pmos 20e-6 1e-6
mn1 2 3 0 0 nmos 10e-6 1e-6
vg 3 0 3
