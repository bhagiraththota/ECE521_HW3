vdd 1 0 5
r1 1 2 1000
m1 2 1 4 0 nmos 10e-6 1e-6
m2 4 3 0 0 nmos 10e-6 1e-6
vg 3 0 3
