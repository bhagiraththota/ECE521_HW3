vcc 1 0 5
r1 1 2 1000
q1 2 3 0 npn
vb 3 0 0.78
