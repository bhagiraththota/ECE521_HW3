m1 3 10 2 2 pmos 150e-6 3e-6
m2 4 11 2 2 pmos 150e-6 3e-6
m3 3 3 101 101 nmos 75e-6 3e-6
m4 4 3 101 101 nmos 75e-6 3e-6
m5 2 1 100 100 pmos 150e-6 3e-6
m6 10 4 101 101 nmos 150e-6 3e-6
m7 10 1 100 100 pmos 150e-6 3e-6
m8 1 1 100 100 pmos 75e-6 3e-6
Iref 1 101 50e-6
vdd 100 0 2.5
vss 101 0 -2.5
vin 11 0 0
